module Lab2(a,b);

	input [0 : 3] a;
	
	output [0 : 6] b;

	assign b[0] = ~((~a[0] & ~a[1] & a[2] & ~a[3]) | (~a[0] & ~a[1] & a[2] & a[3]) | (~a[0] & a[1] & ~a[2] & a[3]) | (~a[0] & a[1] & a[2] & ~a[3]) | (~a[0] & a[1] & a[2] & a[3]) | (a[0] & ~a[1] & ~a[2] & ~a[3]) | (a[0] & ~a[1] & ~a[2] & a[3]) | (a[0] & ~a[1] & a[2] & ~a[3]) | (a[0] & a[1] & ~a[2] & ~a[3]) | (a[0] & a[1] & a[2] & ~a[3]) | (a[0] & a[1] & a[2] & a[3]));
	assign b[1] = ~((~a[0] & ~a[1] & ~a[2] & a[3]) | (~a[0] & ~a[1] & a[2] & ~a[3]) | (~a[0] & ~a[1] & a[2] & a[3]) | (~a[0] & a[1] & ~a[2] & ~a[3]) | (~a[0] & a[1] & a[2] & a[3]) | (a[0] & ~a[1] & ~a[2] & ~a[3]) | (a[0] & ~a[1] & ~a[2] & a[3]) | (a[0] & ~a[1] & a[2] & ~a[3]) | (a[0] & a[1] & ~a[2] & a[3]));
	assign b[2] = ~((~a[0] & ~a[1] & ~a[2] & a[3]) | (~a[0] & ~a[1] & a[2] & a[3]) | (~a[0] & a[1] & ~a[2] & ~a[3]) | (~a[0] & a[1] & ~a[2] & a[3]) | (~a[0] & a[1] & a[2] & ~a[3]) | (~a[0] & a[1] & a[2] & a[3]) | (a[0] & ~a[1] & ~a[2] & ~a[3]) | (a[0] & ~a[1] & ~a[2] & a[3]) | (a[0] & ~a[1] & a[2] & ~a[3]) | (a[0] & ~a[1] & a[2] & a[3]) | (a[0] & a[1] & ~a[2] & a[3]));
	assign b[3] = ~((~a[0] & ~a[1] & a[2] & ~a[3]) | (~a[0] & ~a[1] & a[2] & a[3]) | (~a[0] & a[1] & ~a[2] & a[3]) | (~a[0] & a[1] & a[2] & ~a[3]) | (a[0] & ~a[1] & ~a[2] & ~a[3]) | (a[0] & ~a[1] & ~a[2] & a[3]) | (a[0] & ~a[1] & a[2] & a[3]) | (a[0] & a[1] & ~a[2] & ~a[3]) | (a[0] & a[1] & ~a[2] & a[3]) | (a[0] & a[1] & a[2] & ~a[3]));
	assign b[4] = ~((~a[0] & ~a[1] & a[2] & ~a[3]) | (~a[0] & a[1] & a[2] & ~a[3]) | (a[0] & ~a[1] & ~a[2] & ~a[3]) | (a[0] & ~a[1] & a[2] & ~a[3]) | (a[0] & ~a[1] & a[2] & a[3]) | (a[0] & a[1] & ~a[2] & ~a[3]) | (a[0] & a[1] & ~a[2] & a[3]) | (a[0] & a[1] & a[2] & ~a[3]) | (a[0] & a[1] & a[2] & a[3]));
	
// Equation Reduction for b[5] in minterm form:
// Original expression: (~a[0]~a[1]~a[2]a[3]) + (~a[1]~a[1]a[2]~a[3]) + (~a[0]~a[1]a[2]a[3]) + (~a[0]a[1]a[2]a[3]) + (a[0]a[1]~a[2]a[3]);  
// These are the combinations that give 0 (Which represents LED On in this case)
// 						 	 = (~a[0]~a[1])(~a[2]a[3] + a[2]~a[3] + a[2]a[3]) + (~a[0]a[1]a[2]a[3]) + (a[0]a[1]~a[2]a[3])
// The Expression (~a[2]a[3] + a[2]~a[3] + a[2]a[3]) Will always amount to true in our case because
// (1 & 1) = 1 , (1 & 0) = 1 , (0 & 1) = 1 , (0 & 0) = 0 but this is not necessary in our case becuase it would make a binary value of 0000 which displays nothing
// So, 						 = (~a[0]~a[1])(1) + (~a[0]a[1]a[2]a[3]) + (a[0]a[1]~a[2]a[3])
//      						 = (~a[0]~a[1]) + (~a[0]a[1]a[2]a[3]) + (a[0]a[1]~a[2]a[3])
// And we have reduced the expression

	assign b[5] = (~a[0] & ~a[1]) | (~a[0] & a[1] & a[2] & a[3]) | (a[0] & a[1] & ~a[2] & a[3]);
	
	assign b[6] = ~((~a[0] & ~a[1] & a[2] & ~a[3]) | (~a[0] & ~a[1] & a[2] & a[3]) | (~a[0] & a[1] & ~a[2] & ~a[3]) | (~a[0] & a[1] & ~a[2] & a[3]) | (~a[0] & a[1] & a[2] & ~a[3]) | (a[0] & ~a[1] & ~a[2] & ~a[3]) | (a[0] & ~a[1] & ~a[2] & a[3]) | (a[0] & ~a[1] & a[2] & ~a[3]) | (a[0] & ~a[1] & a[2] & a[3]) | (a[0] & a[1] & ~a[2] & a[3])| (a[0] & a[1] & a[2] & ~a[3]) | (a[0] & a[1] & a[2] & a[3]));

	
endmodule